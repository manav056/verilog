//Interface for verifying dff module

interface dff_if(input bit clk);
    
    logic din;
    logic dout;

endinterface