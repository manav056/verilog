$date
	Sat Sep 14 16:48:26 2024
$end
$version
	Icarus Verilog
$end
$timescale
	1s
$end
$scope module adder8bit_tb $end
$var wire 8 ! out [7:0] $end
$var wire 1 " cout $end
$var reg 8 # a [7:0] $end
$var reg 8 $ b [7:0] $end
$var reg 1 % cin $end
$scope module DUT $end
$var wire 8 & a [7:0] $end
$var wire 8 ' b [7:0] $end
$var wire 1 % cin $end
$var wire 8 ( out [7:0] $end
$var wire 1 " cout $end
$var wire 9 ) carry [8:0] $end
$var parameter 32 * n $end
$scope begin genblk1[0] $end
$var parameter 2 + i $end
$scope module FA0 $end
$var wire 1 , cin $end
$var wire 1 - cout $end
$var wire 1 . sum $end
$var wire 1 / x $end
$var wire 1 0 y $end
$upscope $end
$upscope $end
$scope begin genblk1[1] $end
$var parameter 2 1 i $end
$scope module FA0 $end
$var wire 1 2 cin $end
$var wire 1 3 cout $end
$var wire 1 4 sum $end
$var wire 1 5 x $end
$var wire 1 6 y $end
$upscope $end
$upscope $end
$scope begin genblk1[2] $end
$var parameter 3 7 i $end
$scope module FA0 $end
$var wire 1 8 cin $end
$var wire 1 9 cout $end
$var wire 1 : sum $end
$var wire 1 ; x $end
$var wire 1 < y $end
$upscope $end
$upscope $end
$scope begin genblk1[3] $end
$var parameter 3 = i $end
$scope module FA0 $end
$var wire 1 > cin $end
$var wire 1 ? cout $end
$var wire 1 @ sum $end
$var wire 1 A x $end
$var wire 1 B y $end
$upscope $end
$upscope $end
$scope begin genblk1[4] $end
$var parameter 4 C i $end
$scope module FA0 $end
$var wire 1 D cin $end
$var wire 1 E cout $end
$var wire 1 F sum $end
$var wire 1 G x $end
$var wire 1 H y $end
$upscope $end
$upscope $end
$scope begin genblk1[5] $end
$var parameter 4 I i $end
$scope module FA0 $end
$var wire 1 J cin $end
$var wire 1 K cout $end
$var wire 1 L sum $end
$var wire 1 M x $end
$var wire 1 N y $end
$upscope $end
$upscope $end
$scope begin genblk1[6] $end
$var parameter 4 O i $end
$scope module FA0 $end
$var wire 1 P cin $end
$var wire 1 Q cout $end
$var wire 1 R sum $end
$var wire 1 S x $end
$var wire 1 T y $end
$upscope $end
$upscope $end
$scope begin genblk1[7] $end
$var parameter 4 U i $end
$scope module FA0 $end
$var wire 1 V cin $end
$var wire 1 W cout $end
$var wire 1 X sum $end
$var wire 1 Y x $end
$var wire 1 Z y $end
$upscope $end
$upscope $end
$upscope $end
$upscope $end
$enddefinitions $end
$comment Show the parameter values. $end
$dumpall
b111 U
b110 O
b101 I
b100 C
b11 =
b10 7
b1 1
b0 +
b1000 *
$end
#0
$dumpvars
xZ
xY
xX
xW
xV
xT
xS
xR
xQ
xP
xN
xM
xL
xK
xJ
xH
xG
xF
xE
xD
xB
xA
x@
x?
x>
x<
x;
x:
x9
x8
x6
x5
x4
x3
x2
x0
x/
x.
x-
x,
bx )
bx (
bx '
bx &
x%
bx $
bx #
x"
bx !
$end
#5
0:
0@
0F
0L
0R
0X
14
08
0>
0D
0J
0P
0V
0"
12
03
09
0?
0E
0K
0Q
0W
1-
b10 !
b10 (
0.
0,
10
06
0<
0B
0H
0N
0T
0Z
1/
05
0;
0A
0G
0M
0S
0Y
b10 )
0%
b1 $
b1 '
b1 #
b1 &
#15
b11 !
b11 (
1.
1,
b11 )
1%
#30
b1011 !
b1011 (
1@
1>
1"
19
b100001011 )
1W
1<
1Z
1;
1Y
b10000101 $
b10000101 '
b10000101 #
b10000101 &
